`timescale 1ns / 1ps

module multiplier(product, input1, input2);
	output [7:0] product;
	input [3:0] input1;
	input [3:0] input2;
	
endmodule
